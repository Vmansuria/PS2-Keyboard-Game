-- This project is a game which is implemented for Basys3 using VHDL language for learning purposes.
--It takes inputs from buttons(for game control) and switch(reset) on Basys3, outputs the data on Seven Segment
--Display and on a Monitor that supports VGA standart.

--User controls an object which moves vertically and some bars come in horizontal direction. User tries object to
--avoid from these bars using the up and down buttons on Basys 3. Once one the buttons are pressed the object moves
--in the direction of up/down with constant velocity. Object doesn't stop so user must actively controll it. As the
--time passes, score of the user increase. When the object hits one of the bars or the object hits the uppermost or
--lowermost parts of the screen, game is over and a text indicating this shows up on monitor. At the same time,
--score stop to increase so that user can see their scores.

--It uses 4 modules, one for VGA control, one or Button Debouncer, one for seven segment display on Basys 3, and
--one for the top module which also has the game mechanics.


--This is the top module for the game "Don't Hit The Bars". It has all other modules in it and has the mechanis
--like collision, motion, adjusting the score of the game.

--* vga.vhd and debounce.vhd modules are  taken from VGA project for Basys3 from the user Dries007
--via github. Original codes can be found on https://github.com/dries007/Basys3/tree/master/VGA which
--is licensed under The MIT License (MIT)

--* Two functions draw_char and draw_string are also taken from taken from VGA project for Basys3 from 
--the user Dries007 via github. Those functions are used for demo in that project. Original codes can 
--be found on https://github.com/dries007/Basys3/tree/master/VGA which is licensed 
--under The MIT License (MIT)

--* SevSeg_4digit module is written in SystemVerilog and taken from
--https://dl.dropboxusercontent.com/u/11084576/CS223/SevSeg_4digit.sv which is used in the Bilkent 
--CS 223 course labs and projects.

--Note For the failing timing requirements:
--Timing requirement is not met after the use of code for drawing strings on vga monitor since critical path
--for it is quite long and I didn't want to slow down the clock. However, the program works well because of
--the fact that the text "Game Over!" is displayed at the end of a game and it is centered so it is enough 
--for the purpose. But for further modification, this problem might be attended to.

--Copyright (C) 2017 M. Ali Semi YENIMOL

--Licensed under the TAPR Open Hardware License (www.tapr.org/OHL)

library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.STD_LOGIC_ARITH.ALL;
use IEEE.std_logic_unsigned.all;


entity game is
    Port ( 
        clk : in STD_LOGIC;
        vgaRed : out STD_LOGIC_VECTOR(3 downto 0);
        vgaBlue : out STD_LOGIC_VECTOR(3 downto 0);
        vgaGreen : out STD_LOGIC_VECTOR(3 downto 0);
        Hsync : out STD_LOGIC;
        Vsync : out STD_LOGIC;
--        btnU : in STD_LOGIC;
--        btnD : in STD_LOGIC;
        speed_sw : in STD_LOGIC_VECTOR(2 downto 0);
        reset : in STD_LOGIC;
        seg : out STD_LOGIC_VECTOR(6 downto 0);
        dp : out STD_LOGIC; --For seven segment display on Basys 3
        an : out STD_LOGIC_VECTOR(3 downto 0); --For seven segment display on Basys 3
        ps2c_in : in STD_LOGIC;
        ps2d_in : in STD_LOGIC
    );
end game;

architecture Behavioral of game is
    component Sequential_7Segments_Decoder is
    Port ( 
		
		value : in std_logic_vector(15 downto 0);
		RESET: in std_logic;
		clk : in std_logic;
		dp : out std_logic;
		-- The anodes will be treated as if they are different 
		-- communication channels, which are getting activated and deactivated according to the internal subclock (Sclk)
		channels : out std_logic_vector(3 downto 0);
	    segs : out std_logic_vector(6 downto 0));
    end component;
    
    component ps2keyboard is
        port (resetn, clock: in std_logic;
                ps2c, ps2d: in std_logic;
                DOUT: inout std_logic_vector (8 downto 0);
                code: out std_logic_vector (15 downto 0)
               );
    end component;
    
    signal btn_cnt : natural range 0 to 1000000;
    signal clk_cnt : natural range 0 to 500000;
    
    --All coordinates determines the left corner of an object
    signal posX : natural range 0 to 1280; --x position of the guy
    signal posY : natural range 0 to 1024; --y position of the guy
    
    signal X : natural range 0 to 1280;
    signal Y : natural range 0 to 1024;
    signal Red : natural range 0 to 15;
    signal Green : natural range 0 to 15;
    signal Blue : natural range 0 to 15;
	
	constant sizeOfGuy: natural := 50;
	constant centerX: natural := 640;
	constant centerY: natural := 512;
	constant heightOfBar: natural := 30;
	
	signal moveUp: std_logic; --determines if the guy is moving to up or not
	signal moveDown: std_logic; --determines if the guy is moving to down or not
	signal gameOver: std_logic; --a flag to end up the game
	signal speedOfGuy: natural;
	signal speedOfBars: natural;
	
	--Basically, there might be at most 5 bars can be seen on screen so the lenghts of each bar are
	--also 256 ( 1280/5 = 256)
    type int_array_Y is array (0 to 4) of natural range 0 to 1024;
	type int_array_X is array (0 to 4) of integer range -1280 to 3280;-- Up to 3280 For overflow issues
	type int_array_L is array (0 to 4) of integer range 0 to 500;
	
	--Upcoming bars are storaged as ROM to have a control on the places of bars. But for further
	--modification, random generators might be used as well.
	type int_array_Y_levels is array (0 to 99) of natural range 0 to 1024; 
	type int_array_L_levels is array (0 to 99) of integer range 0 to 300;
	
	--For now, just 2 bars paralel to each other is used. 3 or more bars might be used to increase difficulty
	signal upBarYPositions : int_array_Y;
	signal upBarLengths : int_array_L; --Parallel array with upBarYPositions
	signal upBarXPositions : int_array_X; --Parallel array with upBarYPositions
	
	signal downBarYPositions : int_array_Y;
	signal downBarLengths : int_array_L;
	signal downBarXPositions : int_array_X;
	
	--For later intermediary bars might be needed
	signal currentUpEdge: natural range 0 to 1024 := 0;
	signal currentDownEdge: natural range 0 to 1024 := 0;
	signal frame_count : natural range 0 to 1000000;

	--For next bars as the game progress, used as Rom but random generator implementation might be used as well
	constant upBarYPositionsNext : int_array_Y_levels   := (264,126,170,278,381,376,238,382,282,246,117,345,271,86,369,210,205,318,182,360,52,387,154,168,48,77,254,184,15,206,372,7,79,282,93,264,15,92,12,130,212,66,45,261,170,396,210,135,151,64,11,147,34,217,115,77,258,12,164,204,95,59,76,345,58,29,260,75,330,68,397,130,169,94,43,270,283,195,54,167,347,320,179,88,384,358,220,336,56,334,27,370,383,345,392,6,44,171,280,26);
	constant upBarLengthsNext : int_array_L_levels      := (256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256);	
	constant downBarYPositionsNext : int_array_Y_levels := (550,580,610,640,640,700,700,850,728,697,758,519,831,672,823,530,852,645,697,879,565,589,972,825,927,644,553,792,895,727,1005,605,760,617,791,608,608,794,932,655,670,799,650,892,919,972,550,509,832,548,618,693,884,707,586,653,830,892,656,909,935,871,656,871,889,865,759,636,749,519,729,753,611,850,813,958,879,783,543,999,963,757,734,659,777,529,594,866,512,516,950,686,502,886,912,886,783,872,978,699);
    constant downBarLengthsNext: int_array_L_levels     := (256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256);
    signal indexUpBarNext: natural range 0 to 99;
    signal indexDownBarNext : natural range 0 to 99;
    signal curUp_cnt: natural range 0 to 1000; --curUp_cnt and curDown_cnt are counters for the process where 
    signal curDown_cnt: natural range 0 to 1000;--current edge is determined. They are needed to decrease the frequency of the process
    
    signal in0, in1, in2, in3 : std_logic_vector( 3 downto 0); --Scores given as parameters to sevSeg_4digit
    signal score: natural range 0 to 9999;
    signal score_cnt: natural range 0 to 10000000;
    
    signal Dout : std_logic_vector(8 downto 0) := "000000000";
    signal code_out : std_logic_vector(15 downto 0);
    
--    The MIT License (MIT)
    
--    Copyright (c) 2016 Dries007
    
--    Permission is hereby granted, free of charge, to any person obtaining a copy
--    of this software and associated documentation files (the "Software"), to deal
--    in the Software without restriction, including without limitation the rights
--    to use, copy, modify, merge, publish, distribute, sublicense, and/or sell
--    copies of the Software, and to permit persons to whom the Software is
--    furnished to do so, subject to the following conditions:
    
--    The above copyright notice and this permission notice shall be included in all
--    copies or substantial portions of the Software.
    
--    THE SOFTWARE IS PROVIDED "AS IS", WITHOUT WARRANTY OF ANY KIND, EXPRESS OR
--    IMPLIED, INCLUDING BUT NOT LIMITED TO THE WARRANTIES OF MERCHANTABILITY,
--    FITNESS FOR A PARTICULAR PURPOSE AND NONINFRINGEMENT. IN NO EVENT SHALL THE
--    AUTHORS OR COPYRIGHT HOLDERS BE LIABLE FOR ANY CLAIM, DAMAGES OR OTHER
--    LIABILITY, WHETHER IN AN ACTION OF CONTRACT, TORT OR OTHERWISE, ARISING FROM,
--    OUT OF OR IN CONNECTION WITH THE SOFTWARE OR THE USE OR OTHER DEALINGS IN THE
--    SOFTWARE.
    
    function draw_char(X : natural; Y : natural; char : character) return boolean is
            constant ADDR_WIDTH: integer:=11;
            constant DATA_WIDTH: integer:=8;
            type rom_type is array (0 to 2**ADDR_WIDTH-1) of std_logic_vector(DATA_WIDTH-1 downto 0);
           -- ROM definition
           constant ROM: rom_type:=(   -- 2^11-by-8
           "00000000", -- 0
           "00000000", -- 1
           "00000000", -- 2
           "00000000", -- 3
           "00000000", -- 4
           "00000000", -- 5
           "00000000", -- 6
           "00000000", -- 7
           "00000000", -- 8
           "00000000", -- 9
           "00000000", -- a
           "00000000", -- b
           "00000000", -- c
           "00000000", -- d
           "00000000", -- e
           "00000000", -- f
           -- code x01 ?
           "00000000", -- 0
           "00000000", -- 1
           "01111110", -- 2  ******
           "10000001", -- 3 *      *
           "10100101", -- 4 * *  * *
           "10000001", -- 5 *      *
           "10000001", -- 6 *      *
           "10111101", -- 7 * **** *
           "10011001", -- 8 *  **  *
           "10000001", -- 9 *      *
           "10000001", -- a *      *
           "01111110", -- b  ******
           "00000000", -- c
           "00000000", -- d
           "00000000", -- e
           "00000000", -- f
           -- code x02 ?
           "00000000", -- 0
           "00000000", -- 1
           "01111110", -- 2  ******
           "11111111", -- 3 ********
           "11011011", -- 4 ** ** **
           "11111111", -- 5 ********
           "11111111", -- 6 ********
           "11000011", -- 7 **    **
           "11100111", -- 8 ***  ***
           "11111111", -- 9 ********
           "11111111", -- a ********
           "01111110", -- b  ******
           "00000000", -- c
           "00000000", -- d
           "00000000", -- e
           "00000000", -- f
           -- code x03 ?
           "00000000", -- 0
           "00000000", -- 1
           "00000000", -- 2
           "00000000", -- 3
           "01101100", -- 4  ** **
           "11111110", -- 5 *******
           "11111110", -- 6 *******
           "11111110", -- 7 *******
           "11111110", -- 8 *******
           "01111100", -- 9  *****
           "00111000", -- a   ***
           "00010000", -- b    *
           "00000000", -- c
           "00000000", -- d
           "00000000", -- e
           "00000000", -- f
           -- code x04 ?
           "00000000", -- 0
           "00000000", -- 1
           "00000000", -- 2
           "00000000", -- 3
           "00010000", -- 4    *
           "00111000", -- 5   ***
           "01111100", -- 6  *****
           "11111110", -- 7 *******
           "01111100", -- 8  *****
           "00111000", -- 9   ***
           "00010000", -- a    *
           "00000000", -- b
           "00000000", -- c
           "00000000", -- d
           "00000000", -- e
           "00000000", -- f
           -- code x05 ?
           "00000000", -- 0
           "00000000", -- 1
           "00000000", -- 2
           "00011000", -- 3    **
           "00111100", -- 4   ****
           "00111100", -- 5   ****
           "11100111", -- 6 ***  ***
           "11100111", -- 7 ***  ***
           "11100111", -- 8 ***  ***
           "00011000", -- 9    **
           "00011000", -- a    **
           "00111100", -- b   ****
           "00000000", -- c
           "00000000", -- d
           "00000000", -- e
           "00000000", -- f
           -- code x06 ?
           "00000000", -- 0
           "00000000", -- 1
           "00000000", -- 2
           "00011000", -- 3    **
           "00111100", -- 4   ****
           "01111110", -- 5  ******
           "11111111", -- 6 ********
           "11111111", -- 7 ********
           "01111110", -- 8  ******
           "00011000", -- 9    **
           "00011000", -- a    **
           "00111100", -- b   ****
           "00000000", -- c
           "00000000", -- d
           "00000000", -- e
           "00000000", -- f
           -- code x07 �
           "00000000", -- 0
           "00000000", -- 1
           "00000000", -- 2
           "00000000", -- 3
           "00000000", -- 4
           "00000000", -- 5
           "00011000", -- 6    **
           "00111100", -- 7   ****
           "00111100", -- 8   ****
           "00011000", -- 9    **
           "00000000", -- a
           "00000000", -- b
           "00000000", -- c
           "00000000", -- d
           "00000000", -- e
           "00000000", -- f
           -- code x08 ?
           "11111111", -- 0 ********
           "11111111", -- 1 ********
           "11111111", -- 2 ********
           "11111111", -- 3 ********
           "11111111", -- 4 ********
           "11111111", -- 5 ********
           "11100111", -- 6 ***  ***
           "11000011", -- 7 **    **
           "11000011", -- 8 **    **
           "11100111", -- 9 ***  ***
           "11111111", -- a ********
           "11111111", -- b ********
           "11111111", -- c ********
           "11111111", -- d ********
           "11111111", -- e ********
           "11111111", -- f ********
           -- code x09 ?
           "00000000", -- 0
           "00000000", -- 1
           "00000000", -- 2
           "00000000", -- 3
           "00000000", -- 4
           "00111100", -- 5   ****
           "01100110", -- 6  **  **
           "01000010", -- 7  *    *
           "01000010", -- 8  *    *
           "01100110", -- 9  **  **
           "00111100", -- a   ****
           "00000000", -- b
           "00000000", -- c
           "00000000", -- d
           "00000000", -- e
           "00000000", -- f
           -- code x0a ?
           "11111111", -- 0 ********
           "11111111", -- 1 ********
           "11111111", -- 2 ********
           "11111111", -- 3 ********
           "11111111", -- 4 ********
           "11000011", -- 5 **    **
           "10011001", -- 6 *  **  *
           "10111101", -- 7 * **** *
           "10111101", -- 8 * **** *
           "10011001", -- 9 *  **  *
           "11000011", -- a **    **
           "11111111", -- b ********
           "11111111", -- c ********
           "11111111", -- d ********
           "11111111", -- e ********
           "11111111", -- f ********
           -- code x0b ?
           "00000000", -- 0
           "00000000", -- 1
           "00011110", -- 2    ****
           "00001110", -- 3     ***
           "00011010", -- 4    ** *
           "00110010", -- 5   **  *
           "01111000", -- 6  ****
           "11001100", -- 7 **  **
           "11001100", -- 8 **  **
           "11001100", -- 9 **  **
           "11001100", -- a **  **
           "01111000", -- b  ****
           "00000000", -- c
           "00000000", -- d
           "00000000", -- e
           "00000000", -- f
           -- code x0c ?
           "00000000", -- 0
           "00000000", -- 1
           "00111100", -- 2   ****
           "01100110", -- 3  **  **
           "01100110", -- 4  **  **
           "01100110", -- 5  **  **
           "01100110", -- 6  **  **
           "00111100", -- 7   ****
           "00011000", -- 8    **
           "01111110", -- 9  ******
           "00011000", -- a    **
           "00011000", -- b    **
           "00000000", -- c
           "00000000", -- d
           "00000000", -- e
           "00000000", -- f
           -- code x0d ?
           "00000000", -- 0
           "00000000", -- 1
           "00111111", -- 2   ******
           "00110011", -- 3   **  **
           "00111111", -- 4   ******
           "00110000", -- 5   **
           "00110000", -- 6   **
           "00110000", -- 7   **
           "00110000", -- 8   **
           "01110000", -- 9  ***
           "11110000", -- a ****
           "11100000", -- b ***
           "00000000", -- c
           "00000000", -- d
           "00000000", -- e
           "00000000", -- f
           -- code x0e ?
           "00000000", -- 0
           "00000000", -- 1
           "01111111", -- 2  *******
           "01100011", -- 3  **   **
           "01111111", -- 4  *******
           "01100011", -- 5  **   **
           "01100011", -- 6  **   **
           "01100011", -- 7  **   **
           "01100011", -- 8  **   **
           "01100111", -- 9  **  ***
           "11100111", -- a ***  ***
           "11100110", -- b ***  **
           "11000000", -- c **
           "00000000", -- d
           "00000000", -- e
           "00000000", -- f
           -- code x0f ?
           "00000000", -- 0
           "00000000", -- 1
           "00000000", -- 2
           "00011000", -- 3    **
           "00011000", -- 4    **
           "11011011", -- 5 ** ** **
           "00111100", -- 6   ****
           "11100111", -- 7 ***  ***
           "00111100", -- 8   ****
           "11011011", -- 9 ** ** **
           "00011000", -- a    **
           "00011000", -- b    **
           "00000000", -- c
           "00000000", -- d
           "00000000", -- e
           "00000000", -- f
           -- code x10 ?
           "00000000", -- 0
           "10000000", -- 1 *
           "11000000", -- 2 **
           "11100000", -- 3 ***
           "11110000", -- 4 ****
           "11111000", -- 5 *****
           "11111110", -- 6 *******
           "11111000", -- 7 *****
           "11110000", -- 8 ****
           "11100000", -- 9 ***
           "11000000", -- a **
           "10000000", -- b *
           "00000000", -- c
           "00000000", -- d
           "00000000", -- e
           "00000000", -- f
           -- code x11 ?
           "00000000", -- 0
           "00000010", -- 1       *
           "00000110", -- 2      **
           "00001110", -- 3     ***
           "00011110", -- 4    ****
           "00111110", -- 5   *****
           "11111110", -- 6 *******
           "00111110", -- 7   *****
           "00011110", -- 8    ****
           "00001110", -- 9     ***
           "00000110", -- a      **
           "00000010", -- b       *
           "00000000", -- c
           "00000000", -- d
           "00000000", -- e
           "00000000", -- f
           -- code x12 ?
           "00000000", -- 0
           "00000000", -- 1
           "00011000", -- 2    **
           "00111100", -- 3   ****
           "01111110", -- 4  ******
           "00011000", -- 5    **
           "00011000", -- 6    **
           "00011000", -- 7    **
           "01111110", -- 8  ******
           "00111100", -- 9   ****
           "00011000", -- a    **
           "00000000", -- b
           "00000000", -- c
           "00000000", -- d
           "00000000", -- e
           "00000000", -- f
           -- code x13 ?
           "00000000", -- 0
           "00000000", -- 1
           "01100110", -- 2  **  **
           "01100110", -- 3  **  **
           "01100110", -- 4  **  **
           "01100110", -- 5  **  **
           "01100110", -- 6  **  **
           "01100110", -- 7  **  **
           "01100110", -- 8  **  **
           "00000000", -- 9
           "01100110", -- a  **  **
           "01100110", -- b  **  **
           "00000000", -- c
           "00000000", -- d
           "00000000", -- e
           "00000000", -- f
           -- code x14 �
           "00000000", -- 0
           "00000000", -- 1
           "01111111", -- 2  *******
           "11011011", -- 3 ** ** **
           "11011011", -- 4 ** ** **
           "11011011", -- 5 ** ** **
           "01111011", -- 6  **** **
           "00011011", -- 7    ** **
           "00011011", -- 8    ** **
           "00011011", -- 9    ** **
           "00011011", -- a    ** **
           "00011011", -- b    ** **
           "00000000", -- c
           "00000000", -- d
           "00000000", -- e
           "00000000", -- f
           -- code x15 �
           "00000000", -- 0
           "01111100", -- 1  *****
           "11000110", -- 2 **   **
           "01100000", -- 3  **
           "00111000", -- 4   ***
           "01101100", -- 5  ** **
           "11000110", -- 6 **   **
           "11000110", -- 7 **   **
           "01101100", -- 8  ** **
           "00111000", -- 9   ***
           "00001100", -- a     **
           "11000110", -- b **   **
           "01111100", -- c  *****
           "00000000", -- d
           "00000000", -- e
           "00000000", -- f
           -- code x16 ?
           "00000000", -- 0
           "00000000", -- 1
           "00000000", -- 2
           "00000000", -- 3
           "00000000", -- 4
           "00000000", -- 5
           "00000000", -- 6
           "00000000", -- 7
           "11111110", -- 8 *******
           "11111110", -- 9 *******
           "11111110", -- a *******
           "11111110", -- b *******
           "00000000", -- c
           "00000000", -- d
           "00000000", -- e
           "00000000", -- f
           -- code x17 ?
           "00000000", -- 0
           "00000000", -- 1
           "00011000", -- 2    **
           "00111100", -- 3   ****
           "01111110", -- 4  ******
           "00011000", -- 5    **
           "00011000", -- 6    **
           "00011000", -- 7    **
           "01111110", -- 8  ******
           "00111100", -- 9   ****
           "00011000", -- a    **
           "01111110", -- b  ******
           "00110000", -- c
           "00000000", -- d
           "00000000", -- e
           "00000000", -- f
           -- code x18 ?
           "00000000", -- 0
           "00000000", -- 1
           "00011000", -- 2    **
           "00111100", -- 3   ****
           "01111110", -- 4  ******
           "00011000", -- 5    **
           "00011000", -- 6    **
           "00011000", -- 7    **
           "00011000", -- 8    **
           "00011000", -- 9    **
           "00011000", -- a    **
           "00011000", -- b    **
           "00000000", -- c
           "00000000", -- d
           "00000000", -- e
           "00000000", -- f
           -- code x19 ?
           "00000000", -- 0
           "00000000", -- 1
           "00011000", -- 2    **
           "00011000", -- 3    **
           "00011000", -- 4    **
           "00011000", -- 5    **
           "00011000", -- 6    **
           "00011000", -- 7    **
           "00011000", -- 8    **
           "01111110", -- 9  ******
           "00111100", -- a   ****
           "00011000", -- b    **
           "00000000", -- c
           "00000000", -- d
           "00000000", -- e
           "00000000", -- f
           -- code x1a ?
           "00000000", -- 0
           "00000000", -- 1
           "00000000", -- 2
           "00000000", -- 3
           "00000000", -- 4
           "00011000", -- 5    **
           "00001100", -- 6     **
           "11111110", -- 7 *******
           "00001100", -- 8     **
           "00011000", -- 9    **
           "00000000", -- a
           "00000000", -- b
           "00000000", -- c
           "00000000", -- d
           "00000000", -- e
           "00000000", -- f
           -- code x1b ?
           "00000000", -- 0
           "00000000", -- 1
           "00000000", -- 2
           "00000000", -- 3
           "00000000", -- 4
           "00110000", -- 5   **
           "01100000", -- 6  **
           "11111110", -- 7 *******
           "01100000", -- 8  **
           "00110000", -- 9   **
           "00000000", -- a
           "00000000", -- b
           "00000000", -- c
           "00000000", -- d
           "00000000", -- e
           "00000000", -- f
           -- code x1c ?
           "00000000", -- 0
           "00000000", -- 1
           "00000000", -- 2
           "00000000", -- 3
           "00000000", -- 4
           "00000000", -- 5
           "11000000", -- 6 **
           "11000000", -- 7 **
           "11000000", -- 8 **
           "11111110", -- 9 *******
           "00000000", -- a
           "00000000", -- b
           "00000000", -- c
           "00000000", -- d
           "00000000", -- e
           "00000000", -- f
           -- code x1d ?
           "00000000", -- 0
           "00000000", -- 1
           "00000000", -- 2
           "00000000", -- 3
           "00000000", -- 4
           "00100100", -- 5   *  *
           "01100110", -- 6  **  **
           "11111111", -- 7 ********
           "01100110", -- 8  **  **
           "00100100", -- 9   *  *
           "00000000", -- a
           "00000000", -- b
           "00000000", -- c
           "00000000", -- d
           "00000000", -- e
           "00000000", -- f
           -- code x1e ?
           "00000000", -- 0
           "00000000", -- 1
           "00000000", -- 2
           "00000000", -- 3
           "00010000", -- 4    *
           "00111000", -- 5   ***
           "00111000", -- 6   ***
           "01111100", -- 7  *****
           "01111100", -- 8  *****
           "11111110", -- 9 *******
           "11111110", -- a *******
           "00000000", -- b
           "00000000", -- c
           "00000000", -- d
           "00000000", -- e
           "00000000", -- f
           -- code x1f ?
           "00000000", -- 0
           "00000000", -- 1
           "00000000", -- 2
           "00000000", -- 3
           "11111110", -- 4 *******
           "11111110", -- 5 *******
           "01111100", -- 6  *****
           "01111100", -- 7  *****
           "00111000", -- 8   ***
           "00111000", -- 9   ***
           "00010000", -- a    *
           "00000000", -- b
           "00000000", -- c
           "00000000", -- d
           "00000000", -- e
           "00000000", -- f
           -- code x20 ' '
           "00000000", -- 0
           "00000000", -- 1
           "00000000", -- 2
           "00000000", -- 3
           "00000000", -- 4
           "00000000", -- 5
           "00000000", -- 6
           "00000000", -- 7
           "00000000", -- 8
           "00000000", -- 9
           "00000000", -- a
           "00000000", -- b
           "00000000", -- c
           "00000000", -- d
           "00000000", -- e
           "00000000", -- f
           -- code x21 !
           "00000000", -- 0
           "00000000", -- 1
           "00011000", -- 2    **
           "00111100", -- 3   ****
           "00111100", -- 4   ****
           "00111100", -- 5   ****
           "00011000", -- 6    **
           "00011000", -- 7    **
           "00011000", -- 8    **
           "00000000", -- 9
           "00011000", -- a    **
           "00011000", -- b    **
           "00000000", -- c
           "00000000", -- d
           "00000000", -- e
           "00000000", -- f
           -- code x22 "
           "00000000", -- 0
           "01100110", -- 1  **  **
           "01100110", -- 2  **  **
           "01100110", -- 3  **  **
           "00100100", -- 4   *  *
           "00000000", -- 5
           "00000000", -- 6
           "00000000", -- 7
           "00000000", -- 8
           "00000000", -- 9
           "00000000", -- a
           "00000000", -- b
           "00000000", -- c
           "00000000", -- d
           "00000000", -- e
           "00000000", -- f
           -- code x23 #
           "00000000", -- 0
           "00000000", -- 1
           "00000000", -- 2
           "01101100", -- 3  ** **
           "01101100", -- 4  ** **
           "11111110", -- 5 *******
           "01101100", -- 6  ** **
           "01101100", -- 7  ** **
           "01101100", -- 8  ** **
           "11111110", -- 9 *******
           "01101100", -- a  ** **
           "01101100", -- b  ** **
           "00000000", -- c
           "00000000", -- d
           "00000000", -- e
           "00000000", -- f
           -- code x24 $
           "00011000", -- 0     **
           "00011000", -- 1     **
           "01111100", -- 2   *****
           "11000110", -- 3  **   **
           "11000010", -- 4  **    *
           "11000000", -- 5  **
           "01111100", -- 6   *****
           "00000110", -- 7       **
           "00000110", -- 8       **
           "10000110", -- 9  *    **
           "11000110", -- a  **   **
           "01111100", -- b   *****
           "00011000", -- c     **
           "00011000", -- d     **
           "00000000", -- e
           "00000000", -- f
           -- code x25 %
           "00000000", -- 0
           "00000000", -- 1
           "00000000", -- 2
           "00000000", -- 3
           "11000010", -- 4 **    *
           "11000110", -- 5 **   **
           "00001100", -- 6     **
           "00011000", -- 7    **
           "00110000", -- 8   **
           "01100000", -- 9  **
           "11000110", -- a **   **
           "10000110", -- b *    **
           "00000000", -- c
           "00000000", -- d
           "00000000", -- e
           "00000000", -- f
           -- code x26 &
           "00000000", -- 0
           "00000000", -- 1
           "00111000", -- 2   ***
           "01101100", -- 3  ** **
           "01101100", -- 4  ** **
           "00111000", -- 5   ***
           "01110110", -- 6  *** **
           "11011100", -- 7 ** ***
           "11001100", -- 8 **  **
           "11001100", -- 9 **  **
           "11001100", -- a **  **
           "01110110", -- b  *** **
           "00000000", -- c
           "00000000", -- d
           "00000000", -- e
           "00000000", -- f
           -- code x27 '
           "00000000", -- 0
           "00110000", -- 1   **
           "00110000", -- 2   **
           "00110000", -- 3   **
           "01100000", -- 4  **
           "00000000", -- 5
           "00000000", -- 6
           "00000000", -- 7
           "00000000", -- 8
           "00000000", -- 9
           "00000000", -- a
           "00000000", -- b
           "00000000", -- c
           "00000000", -- d
           "00000000", -- e
           "00000000", -- f
           -- code x28 (
           "00000000", -- 0
           "00000000", -- 1
           "00001100", -- 2     **
           "00011000", -- 3    **
           "00110000", -- 4   **
           "00110000", -- 5   **
           "00110000", -- 6   **
           "00110000", -- 7   **
           "00110000", -- 8   **
           "00110000", -- 9   **
           "00011000", -- a    **
           "00001100", -- b     **
           "00000000", -- c
           "00000000", -- d
           "00000000", -- e
           "00000000", -- f
           -- code x29 )
           "00000000", -- 0
           "00000000", -- 1
           "00110000", -- 2   **
           "00011000", -- 3    **
           "00001100", -- 4     **
           "00001100", -- 5     **
           "00001100", -- 6     **
           "00001100", -- 7     **
           "00001100", -- 8     **
           "00001100", -- 9     **
           "00011000", -- a    **
           "00110000", -- b   **
           "00000000", -- c
           "00000000", -- d
           "00000000", -- e
           "00000000", -- f
           -- code x2a *
           "00000000", -- 0
           "00000000", -- 1
           "00000000", -- 2
           "00000000", -- 3
           "00000000", -- 4
           "01100110", -- 5  **  **
           "00111100", -- 6   ****
           "11111111", -- 7 ********
           "00111100", -- 8   ****
           "01100110", -- 9  **  **
           "00000000", -- a
           "00000000", -- b
           "00000000", -- c
           "00000000", -- d
           "00000000", -- e
           "00000000", -- f
           -- code x2b +
           "00000000", -- 0
           "00000000", -- 1
           "00000000", -- 2
           "00000000", -- 3
           "00000000", -- 4
           "00011000", -- 5    **
           "00011000", -- 6    **
           "01111110", -- 7  ******
           "00011000", -- 8    **
           "00011000", -- 9    **
           "00000000", -- a
           "00000000", -- b
           "00000000", -- c
           "00000000", -- d
           "00000000", -- e
           "00000000", -- f
           -- code x2c ,
           "00000000", -- 0
           "00000000", -- 1
           "00000000", -- 2
           "00000000", -- 3
           "00000000", -- 4
           "00000000", -- 5
           "00000000", -- 6
           "00000000", -- 7
           "00000000", -- 8
           "00011000", -- 9    **
           "00011000", -- a    **
           "00011000", -- b    **
           "00110000", -- c   **
           "00000000", -- d
           "00000000", -- e
           "00000000", -- f
           -- code x2d -
           "00000000", -- 0
           "00000000", -- 1
           "00000000", -- 2
           "00000000", -- 3
           "00000000", -- 4
           "00000000", -- 5
           "00000000", -- 6
           "01111110", -- 7  ******
           "00000000", -- 8
           "00000000", -- 9
           "00000000", -- a
           "00000000", -- b
           "00000000", -- c
           "00000000", -- d
           "00000000", -- e
           "00000000", -- f
           -- code x2e  .
           "00000000", -- 0
           "00000000", -- 1
           "00000000", -- 2
           "00000000", -- 3
           "00000000", -- 4
           "00000000", -- 5
           "00000000", -- 6
           "00000000", -- 7
           "00000000", -- 8
           "00000000", -- 9
           "00011000", -- a    **
           "00011000", -- b    **
           "00000000", -- c
           "00000000", -- d
           "00000000", -- e
           "00000000", -- f
           -- code x2f /
           "00000000", -- 0
           "00000000", -- 1
           "00000000", -- 2
           "00000000", -- 3
           "00000010", -- 4       *
           "00000110", -- 5      **
           "00001100", -- 6     **
           "00011000", -- 7    **
           "00110000", -- 8   **
           "01100000", -- 9  **
           "11000000", -- a **
           "10000000", -- b *
           "00000000", -- c
           "00000000", -- d
           "00000000", -- e
           "00000000", -- f
           -- code x30
           "00000000", -- 0
           "00000000", -- 1
           "01111100", -- 2  *****
           "11000110", -- 3 **   **
           "11000110", -- 4 **   **
           "11001110", -- 5 **  ***
           "11011110", -- 6 ** ****
           "11110110", -- 7 **** **
           "11100110", -- 8 ***  **
           "11000110", -- 9 **   **
           "11000110", -- a **   **
           "01111100", -- b  *****
           "00000000", -- c
           "00000000", -- d
           "00000000", -- e
           "00000000", -- f
           -- code x31 
           "00000000", -- 0
           "00000000", -- 1
           "00011000", -- 2
           "00111000", -- 3
           "01111000", -- 4    **
           "00011000", -- 5   ***
           "00011000", -- 6  ****
           "00011000", -- 7    **
           "00011000", -- 8    **
           "00011000", -- 9    **
           "00011000", -- a    **
           "01111110", -- b    **
           "00000000", -- c    **
           "00000000", -- d  ******
           "00000000", -- e
           "00000000", -- f
           -- code x32
           "00000000", -- 0
           "00000000", -- 1
           "01111100", -- 2  *****
           "11000110", -- 3 **   **
           "00000110", -- 4      **
           "00001100", -- 5     **
           "00011000", -- 6    **
           "00110000", -- 7   **
           "01100000", -- 8  **
           "11000000", -- 9 **
           "11000110", -- a **   **
           "11111110", -- b *******
           "00000000", -- c
           "00000000", -- d
           "00000000", -- e
           "00000000", -- f
           -- code x33
           "00000000", -- 0
           "00000000", -- 1
           "01111100", -- 2  *****
           "11000110", -- 3 **   **
           "00000110", -- 4      **
           "00000110", -- 5      **
           "00111100", -- 6   ****
           "00000110", -- 7      **
           "00000110", -- 8      **
           "00000110", -- 9      **
           "11000110", -- a **   **
           "01111100", -- b  *****
           "00000000", -- c
           "00000000", -- d
           "00000000", -- e
           "00000000", -- f
           -- code x34
           "00000000", -- 0
           "00000000", -- 1
           "00001100", -- 2     **
           "00011100", -- 3    ***
           "00111100", -- 4   ****
           "01101100", -- 5  ** **
           "11001100", -- 6 **  **
           "11111110", -- 7 *******
           "00001100", -- 8     **
           "00001100", -- 9     **
           "00001100", -- a     **
           "00011110", -- b    ****
           "00000000", -- c
           "00000000", -- d
           "00000000", -- e
           "00000000", -- f
           -- code x35
           "00000000", -- 0
           "00000000", -- 1
           "11111110", -- 2 *******
           "11000000", -- 3 **
           "11000000", -- 4 **
           "11000000", -- 5 **
           "11111100", -- 6 ******
           "00000110", -- 7      **
           "00000110", -- 8      **
           "00000110", -- 9      **
           "11000110", -- a **   **
           "01111100", -- b  *****
           "00000000", -- c
           "00000000", -- d
           "00000000", -- e
           "00000000", -- f
           -- code x36
           "00000000", -- 0
           "00000000", -- 1
           "00111000", -- 2   ***
           "01100000", -- 3  **
           "11000000", -- 4 **
           "11000000", -- 5 **
           "11111100", -- 6 ******
           "11000110", -- 7 **   **
           "11000110", -- 8 **   **
           "11000110", -- 9 **   **
           "11000110", -- a **   **
           "01111100", -- b  *****
           "00000000", -- c
           "00000000", -- d
           "00000000", -- e
           "00000000", -- f
           -- code x37
           "00000000", -- 0
           "00000000", -- 1
           "11111110", -- 2 *******
           "11000110", -- 3 **   **
           "00000110", -- 4      **
           "00000110", -- 5      **
           "00001100", -- 6     **
           "00011000", -- 7    **
           "00110000", -- 8   **
           "00110000", -- 9   **
           "00110000", -- a   **
           "00110000", -- b   **
           "00000000", -- c
           "00000000", -- d
           "00000000", -- e
           "00000000", -- f
           -- code x38
           "00000000", -- 0
           "00000000", -- 1
           "01111100", -- 2  *****
           "11000110", -- 3 **   **
           "11000110", -- 4 **   **
           "11000110", -- 5 **   **
           "01111100", -- 6  *****
           "11000110", -- 7 **   **
           "11000110", -- 8 **   **
           "11000110", -- 9 **   **
           "11000110", -- a **   **
           "01111100", -- b  *****
           "00000000", -- c
           "00000000", -- d
           "00000000", -- e
           "00000000", -- f
           -- code x39
           "00000000", -- 0
           "00000000", -- 1
           "01111100", -- 2  *****
           "11000110", -- 3 **   **
           "11000110", -- 4 **   **
           "11000110", -- 5 **   **
           "01111110", -- 6  ******
           "00000110", -- 7      **
           "00000110", -- 8      **
           "00000110", -- 9      **
           "00001100", -- a     **
           "01111000", -- b  ****
           "00000000", -- c
           "00000000", -- d
           "00000000", -- e
           "00000000", -- f
           -- code x3a :
           "00000000", -- 0
           "00000000", -- 1
           "00000000", -- 2
           "00000000", -- 3
           "00011000", -- 4    **
           "00011000", -- 5    **
           "00000000", -- 6
           "00000000", -- 7
           "00000000", -- 8
           "00011000", -- 9    **
           "00011000", -- a    **
           "00000000", -- b
           "00000000", -- c
           "00000000", -- d
           "00000000", -- e
           "00000000", -- f
           -- code x3b ;
           "00000000", -- 0
           "00000000", -- 1
           "00000000", -- 2
           "00000000", -- 3
           "00011000", -- 4    **
           "00011000", -- 5    **
           "00000000", -- 6
           "00000000", -- 7
           "00000000", -- 8
           "00011000", -- 9    **
           "00011000", -- a    **
           "00110000", -- b   **
           "00000000", -- c
           "00000000", -- d
           "00000000", -- e
           "00000000", -- f
           -- code x3c <
           "00000000", -- 0
           "00000000", -- 1
           "00000000", -- 2
           "00000110", -- 3      **
           "00001100", -- 4     **
           "00011000", -- 5    **
           "00110000", -- 6   **
           "01100000", -- 7  **
           "00110000", -- 8   **
           "00011000", -- 9    **
           "00001100", -- a     **
           "00000110", -- b      **
           "00000000", -- c
           "00000000", -- d
           "00000000", -- e
           "00000000", -- f
           -- code x3d =
           "00000000", -- 0
           "00000000", -- 1
           "00000000", -- 2
           "00000000", -- 3
           "00000000", -- 4
           "01111110", -- 5  ******
           "00000000", -- 6
           "00000000", -- 7
           "01111110", -- 8  ******
           "00000000", -- 9
           "00000000", -- a
           "00000000", -- b
           "00000000", -- c
           "00000000", -- d
           "00000000", -- e
           "00000000", -- f
           -- code x3e >
           "00000000", -- 0
           "00000000", -- 1
           "00000000", -- 2
           "01100000", -- 3  **
           "00110000", -- 4   **
           "00011000", -- 5    **
           "00001100", -- 6     **
           "00000110", -- 7      **
           "00001100", -- 8     **
           "00011000", -- 9    **
           "00110000", -- a   **
           "01100000", -- b  **
           "00000000", -- c
           "00000000", -- d
           "00000000", -- e
           "00000000", -- f
           -- code x3f ?
           "00000000", -- 0
           "00000000", -- 1
           "01111100", -- 2  *****
           "11000110", -- 3 **   **
           "11000110", -- 4 **   **
           "00001100", -- 5     **
           "00011000", -- 6    **
           "00011000", -- 7    **
           "00011000", -- 8    **
           "00000000", -- 9
           "00011000", -- a    **
           "00011000", -- b    **
           "00000000", -- c
           "00000000", -- d
           "00000000", -- e
           "00000000", -- f
           -- code x40 @
           "00000000", -- 0
           "00000000", -- 1
           "01111100", -- 2  *****
           "11000110", -- 3 **   **
           "11000110", -- 4 **   **
           "11000110", -- 5 **   **
           "11011110", -- 6 ** ****
           "11011110", -- 7 ** ****
           "11011110", -- 8 ** ****
           "11011100", -- 9 ** ***
           "11000000", -- a **
           "01111100", -- b  *****
           "00000000", -- c
           "00000000", -- d
           "00000000", -- e
           "00000000", -- f
           -- code x41
           "00000000", -- 0
           "00000000", -- 1
           "00010000", -- 2    *
           "00111000", -- 3   ***
           "01101100", -- 4  ** **
           "11000110", -- 5 **   **
           "11000110", -- 6 **   **
           "11111110", -- 7 *******
           "11000110", -- 8 **   **
           "11000110", -- 9 **   **
           "11000110", -- a **   **
           "11000110", -- b **   **
           "00000000", -- c
           "00000000", -- d
           "00000000", -- e
           "00000000", -- f
           -- code x42
           "00000000", -- 0
           "00000000", -- 1
           "11111100", -- 2 ******
           "01100110", -- 3  **  **
           "01100110", -- 4  **  **
           "01100110", -- 5  **  **
           "01111100", -- 6  *****
           "01100110", -- 7  **  **
           "01100110", -- 8  **  **
           "01100110", -- 9  **  **
           "01100110", -- a  **  **
           "11111100", -- b ******
           "00000000", -- c
           "00000000", -- d
           "00000000", -- e
           "00000000", -- f
           -- code x43
           "00000000", -- 0
           "00000000", -- 1
           "00111100", -- 2   ****
           "01100110", -- 3  **  **
           "11000010", -- 4 **    *
           "11000000", -- 5 **
           "11000000", -- 6 **
           "11000000", -- 7 **
           "11000000", -- 8 **
           "11000010", -- 9 **    *
           "01100110", -- a  **  **
           "00111100", -- b   ****
           "00000000", -- c
           "00000000", -- d
           "00000000", -- e
           "00000000", -- f
           -- code x44
           "00000000", -- 0
           "00000000", -- 1
           "11111000", -- 2 *****
           "01101100", -- 3  ** **
           "01100110", -- 4  **  **
           "01100110", -- 5  **  **
           "01100110", -- 6  **  **
           "01100110", -- 7  **  **
           "01100110", -- 8  **  **
           "01100110", -- 9  **  **
           "01101100", -- a  ** **
           "11111000", -- b *****
           "00000000", -- c
           "00000000", -- d
           "00000000", -- e
           "00000000", -- f
           -- code x45
           "00000000", -- 0
           "00000000", -- 1
           "11111110", -- 2 *******
           "01100110", -- 3  **  **
           "01100010", -- 4  **   *
           "01101000", -- 5  ** *
           "01111000", -- 6  ****
           "01101000", -- 7  ** *
           "01100000", -- 8  **
           "01100010", -- 9  **   *
           "01100110", -- a  **  **
           "11111110", -- b *******
           "00000000", -- c
           "00000000", -- d
           "00000000", -- e
           "00000000", -- f
           -- code x46
           "00000000", -- 0
           "00000000", -- 1
           "11111110", -- 2 *******
           "01100110", -- 3  **  **
           "01100010", -- 4  **   *
           "01101000", -- 5  ** *
           "01111000", -- 6  ****
           "01101000", -- 7  ** *
           "01100000", -- 8  **
           "01100000", -- 9  **
           "01100000", -- a  **
           "11110000", -- b ****
           "00000000", -- c
           "00000000", -- d
           "00000000", -- e
           "00000000", -- f
           -- code x47
           "00000000", -- 0
           "00000000", -- 1
           "00111100", -- 2   ****
           "01100110", -- 3  **  **
           "11000010", -- 4 **    *
           "11000000", -- 5 **
           "11000000", -- 6 **
           "11011110", -- 7 ** ****
           "11000110", -- 8 **   **
           "11000110", -- 9 **   **
           "01100110", -- a  **  **
           "00111010", -- b   *** *
           "00000000", -- c
           "00000000", -- d
           "00000000", -- e
           "00000000", -- f
           -- code x48
           "00000000", -- 0
           "00000000", -- 1
           "11000110", -- 2 **   **
           "11000110", -- 3 **   **
           "11000110", -- 4 **   **
           "11000110", -- 5 **   **
           "11111110", -- 6 *******
           "11000110", -- 7 **   **
           "11000110", -- 8 **   **
           "11000110", -- 9 **   **
           "11000110", -- a **   **
           "11000110", -- b **   **
           "00000000", -- c
           "00000000", -- d
           "00000000", -- e
           "00000000", -- f
           -- code x49
           "00000000", -- 0
           "00000000", -- 1
           "00111100", -- 2   ****
           "00011000", -- 3    **
           "00011000", -- 4    **
           "00011000", -- 5    **
           "00011000", -- 6    **
           "00011000", -- 7    **
           "00011000", -- 8    **
           "00011000", -- 9    **
           "00011000", -- a    **
           "00111100", -- b   ****
           "00000000", -- c
           "00000000", -- d
           "00000000", -- e
           "00000000", -- f
           -- code x4a
           "00000000", -- 0
           "00000000", -- 1
           "00011110", -- 2    ****
           "00001100", -- 3     **
           "00001100", -- 4     **
           "00001100", -- 5     **
           "00001100", -- 6     **
           "00001100", -- 7     **
           "11001100", -- 8 **  **
           "11001100", -- 9 **  **
           "11001100", -- a **  **
           "01111000", -- b  ****
           "00000000", -- c
           "00000000", -- d
           "00000000", -- e
           "00000000", -- f
           -- code x4b
           "00000000", -- 0
           "00000000", -- 1
           "11100110", -- 2 ***  **
           "01100110", -- 3  **  **
           "01100110", -- 4  **  **
           "01101100", -- 5  ** **
           "01111000", -- 6  ****
           "01111000", -- 7  ****
           "01101100", -- 8  ** **
           "01100110", -- 9  **  **
           "01100110", -- a  **  **
           "11100110", -- b ***  **
           "00000000", -- c
           "00000000", -- d
           "00000000", -- e
           "00000000", -- f
           -- code x4c
           "00000000", -- 0
           "00000000", -- 1
           "11110000", -- 2 ****
           "01100000", -- 3  **
           "01100000", -- 4  **
           "01100000", -- 5  **
           "01100000", -- 6  **
           "01100000", -- 7  **
           "01100000", -- 8  **
           "01100010", -- 9  **   *
           "01100110", -- a  **  **
           "11111110", -- b *******
           "00000000", -- c
           "00000000", -- d
           "00000000", -- e
           "00000000", -- f
           -- code x4d
           "00000000", -- 0
           "00000000", -- 1
           "11000011", -- 2 **    **
           "11100111", -- 3 ***  ***
           "11111111", -- 4 ********
           "11111111", -- 5 ********
           "11011011", -- 6 ** ** **
           "11000011", -- 7 **    **
           "11000011", -- 8 **    **
           "11000011", -- 9 **    **
           "11000011", -- a **    **
           "11000011", -- b **    **
           "00000000", -- c
           "00000000", -- d
           "00000000", -- e
           "00000000", -- f
           -- code x4e
           "00000000", -- 0
           "00000000", -- 1
           "11000110", -- 2 **   **
           "11100110", -- 3 ***  **
           "11110110", -- 4 **** **
           "11111110", -- 5 *******
           "11011110", -- 6 ** ****
           "11001110", -- 7 **  ***
           "11000110", -- 8 **   **
           "11000110", -- 9 **   **
           "11000110", -- a **   **
           "11000110", -- b **   **
           "00000000", -- c
           "00000000", -- d
           "00000000", -- e
           "00000000", -- f
           -- code x4f
           "00000000", -- 0
           "00000000", -- 1
           "01111100", -- 2  *****
           "11000110", -- 3 **   **
           "11000110", -- 4 **   **
           "11000110", -- 5 **   **
           "11000110", -- 6 **   **
           "11000110", -- 7 **   **
           "11000110", -- 8 **   **
           "11000110", -- 9 **   **
           "11000110", -- a **   **
           "01111100", -- b  *****
           "00000000", -- c
           "00000000", -- d
           "00000000", -- e
           "00000000", -- f
           -- code x50
           "00000000", -- 0
           "00000000", -- 1
           "11111100", -- 2 ******
           "01100110", -- 3  **  **
           "01100110", -- 4  **  **
           "01100110", -- 5  **  **
           "01111100", -- 6  *****
           "01100000", -- 7  **
           "01100000", -- 8  **
           "01100000", -- 9  **
           "01100000", -- a  **
           "11110000", -- b ****
           "00000000", -- c
           "00000000", -- d
           "00000000", -- e
           "00000000", -- f
           -- code x510
           "00000000", -- 0
           "00000000", -- 1
           "01111100", -- 2  *****
           "11000110", -- 3 **   **
           "11000110", -- 4 **   **
           "11000110", -- 5 **   **
           "11000110", -- 6 **   **
           "11000110", -- 7 **   **
           "11000110", -- 8 **   **
           "11010110", -- 9 ** * **
           "11011110", -- a ** ****
           "01111100", -- b  *****
           "00001100", -- c     **
           "00001110", -- d     ***
           "00000000", -- e
           "00000000", -- f
           -- code x52
           "00000000", -- 0
           "00000000", -- 1
           "11111100", -- 2 ******
           "01100110", -- 3  **  **
           "01100110", -- 4  **  **
           "01100110", -- 5  **  **
           "01111100", -- 6  *****
           "01101100", -- 7  ** **
           "01100110", -- 8  **  **
           "01100110", -- 9  **  **
           "01100110", -- a  **  **
           "11100110", -- b ***  **
           "00000000", -- c
           "00000000", -- d
           "00000000", -- e
           "00000000", -- f
           -- code x53
           "00000000", -- 0
           "00000000", -- 1
           "01111100", -- 2  *****
           "11000110", -- 3 **   **
           "11000110", -- 4 **   **
           "01100000", -- 5  **
           "00111000", -- 6   ***
           "00001100", -- 7     **
           "00000110", -- 8      **
           "11000110", -- 9 **   **
           "11000110", -- a **   **
           "01111100", -- b  *****
           "00000000", -- c
           "00000000", -- d
           "00000000", -- e
           "00000000", -- f
           -- code x54
           "00000000", -- 0
           "00000000", -- 1
           "11111111", -- 2 ********
           "11011011", -- 3 ** ** **
           "10011001", -- 4 *  **  *
           "00011000", -- 5    **
           "00011000", -- 6    **
           "00011000", -- 7    **
           "00011000", -- 8    **
           "00011000", -- 9    **
           "00011000", -- a    **
           "00111100", -- b   ****
           "00000000", -- c
           "00000000", -- d
           "00000000", -- e
           "00000000", -- f
           -- code x55
           "00000000", -- 0
           "00000000", -- 1
           "11000110", -- 2 **   **
           "11000110", -- 3 **   **
           "11000110", -- 4 **   **
           "11000110", -- 5 **   **
           "11000110", -- 6 **   **
           "11000110", -- 7 **   **
           "11000110", -- 8 **   **
           "11000110", -- 9 **   **
           "11000110", -- a **   **
           "01111100", -- b  *****
           "00000000", -- c
           "00000000", -- d
           "00000000", -- e
           "00000000", -- f
           -- code x56
           "00000000", -- 0
           "00000000", -- 1
           "11000011", -- 2 **    **
           "11000011", -- 3 **    **
           "11000011", -- 4 **    **
           "11000011", -- 5 **    **
           "11000011", -- 6 **    **
           "11000011", -- 7 **    **
           "11000011", -- 8 **    **
           "01100110", -- 9  **  **
           "00111100", -- a   ****
           "00011000", -- b    **
           "00000000", -- c
           "00000000", -- d
           "00000000", -- e
           "00000000", -- f
           -- code x57
           "00000000", -- 0
           "00000000", -- 1
           "11000011", -- 2 **    **
           "11000011", -- 3 **    **
           "11000011", -- 4 **    **
           "11000011", -- 5 **    **
           "11000011", -- 6 **    **
           "11011011", -- 7 ** ** **
           "11011011", -- 8 ** ** **
           "11111111", -- 9 ********
           "01100110", -- a  **  **
           "01100110", -- b  **  **
           "00000000", -- c
           "00000000", -- d
           "00000000", -- e
           "00000000", -- f
        
           -- code x58
           "00000000", -- 0
           "00000000", -- 1
           "11000011", -- 2 **    **
           "11000011", -- 3 **    **
           "01100110", -- 4  **  **
           "00111100", -- 5   ****
           "00011000", -- 6    **
           "00011000", -- 7    **
           "00111100", -- 8   ****
           "01100110", -- 9  **  **
           "11000011", -- a **    **
           "11000011", -- b **    **
           "00000000", -- c
           "00000000", -- d
           "00000000", -- e
           "00000000", -- f
           -- code x59
           "00000000", -- 0
           "00000000", -- 1
           "11000011", -- 2 **    **
           "11000011", -- 3 **    **
           "11000011", -- 4 **    **
           "01100110", -- 5  **  **
           "00111100", -- 6   ****
           "00011000", -- 7    **
           "00011000", -- 8    **
           "00011000", -- 9    **
           "00011000", -- a    **
           "00111100", -- b   ****
           "00000000", -- c
           "00000000", -- d
           "00000000", -- e
           "00000000", -- f
           -- code x5a
           "00000000", -- 0
           "00000000", -- 1
           "11111111", -- 2 ********
           "11000011", -- 3 **    **
           "10000110", -- 4 *    **
           "00001100", -- 5     **
           "00011000", -- 6    **
           "00110000", -- 7   **
           "01100000", -- 8  **
           "11000001", -- 9 **     *
           "11000011", -- a **    **
           "11111111", -- b ********
           "00000000", -- c
           "00000000", -- d
           "00000000", -- e
           "00000000", -- f
           -- code x5b
           "00000000", -- 0
           "00000000", -- 1
           "00111100", -- 2   ****
           "00110000", -- 3   **
           "00110000", -- 4   **
           "00110000", -- 5   **
           "00110000", -- 6   **
           "00110000", -- 7   **
           "00110000", -- 8   **
           "00110000", -- 9   **
           "00110000", -- a   **
           "00111100", -- b   ****
           "00000000", -- c
           "00000000", -- d
           "00000000", -- e
           "00000000", -- f
           -- code x5c
           "00000000", -- 0
           "00000000", -- 1
           "00000000", -- 2
           "10000000", -- 3 *
           "11000000", -- 4 **
           "11100000", -- 5 ***
           "01110000", -- 6  ***
           "00111000", -- 7   ***
           "00011100", -- 8    ***
           "00001110", -- 9     ***
           "00000110", -- a      **
           "00000010", -- b       *
           "00000000", -- c
           "00000000", -- d
           "00000000", -- e
           "00000000", -- f
           -- code x5d
           "00000000", -- 0
           "00000000", -- 1
           "00111100", -- 2   ****
           "00001100", -- 3     **
           "00001100", -- 4     **
           "00001100", -- 5     **
           "00001100", -- 6     **
           "00001100", -- 7     **
           "00001100", -- 8     **
           "00001100", -- 9     **
           "00001100", -- a     **
           "00111100", -- b   ****
           "00000000", -- c
           "00000000", -- d
           "00000000", -- e
           "00000000", -- f
           -- code x5e
           "00010000", -- 0    *
           "00111000", -- 1   ***
           "01101100", -- 2  ** **
           "11000110", -- 3 **   **
           "00000000", -- 4
           "00000000", -- 5
           "00000000", -- 6
           "00000000", -- 7
           "00000000", -- 8
           "00000000", -- 9
           "00000000", -- a
           "00000000", -- b
           "00000000", -- c
           "00000000", -- d
           "00000000", -- e
           "00000000", -- f
           -- code x5f
           "00000000", -- 0
           "00000000", -- 1
           "00000000", -- 2
           "00000000", -- 3
           "00000000", -- 4
           "00000000", -- 5
           "00000000", -- 6
           "00000000", -- 7
           "00000000", -- 8
           "00000000", -- 9
           "00000000", -- a
           "00000000", -- b
           "00000000", -- c
           "11111111", -- d ********
           "00000000", -- e
           "00000000", -- f
           -- code x60
           "00110000", -- 0   **
           "00110000", -- 1   **
           "00011000", -- 2    **
           "00000000", -- 3
           "00000000", -- 4
           "00000000", -- 5
           "00000000", -- 6
           "00000000", -- 7
           "00000000", -- 8
           "00000000", -- 9
           "00000000", -- a
           "00000000", -- b
           "00000000", -- c
           "00000000", -- d
           "00000000", -- e
           "00000000", -- f
           -- code x61
           "00000000", -- 0
           "00000000", -- 1
           "00000000", -- 2
           "00000000", -- 3
           "00000000", -- 4
           "01111000", -- 5  ****
           "00001100", -- 6     **
           "01111100", -- 7  *****
           "11001100", -- 8 **  **
           "11001100", -- 9 **  **
           "11001100", -- a **  **
           "01110110", -- b  *** **
           "00000000", -- c
           "00000000", -- d
           "00000000", -- e
           "00000000", -- f
           -- code x62
           "00000000", -- 0
           "00000000", -- 1
           "11100000", -- 2  ***
           "01100000", -- 3   **
           "01100000", -- 4   **
           "01111000", -- 5   ****
           "01101100", -- 6   ** **
           "01100110", -- 7   **  **
           "01100110", -- 8   **  **
           "01100110", -- 9   **  **
           "01100110", -- a   **  **
           "01111100", -- b   *****
           "00000000", -- c
           "00000000", -- d
           "00000000", -- e
           "00000000", -- f
           -- code x63
           "00000000", -- 0
           "00000000", -- 1
           "00000000", -- 2
           "00000000", -- 3
           "00000000", -- 4
           "01111100", -- 5  *****
           "11000110", -- 6 **   **
           "11000000", -- 7 **
           "11000000", -- 8 **
           "11000000", -- 9 **
           "11000110", -- a **   **
           "01111100", -- b  *****
           "00000000", -- c
           "00000000", -- d
           "00000000", -- e
           "00000000", -- f
           -- code x64
           "00000000", -- 0
           "00000000", -- 1
           "00011100", -- 2    ***
           "00001100", -- 3     **
           "00001100", -- 4     **
           "00111100", -- 5   ****
           "01101100", -- 6  ** **
           "11001100", -- 7 **  **
           "11001100", -- 8 **  **
           "11001100", -- 9 **  **
           "11001100", -- a **  **
           "01110110", -- b  *** **
           "00000000", -- c
           "00000000", -- d
           "00000000", -- e
           "00000000", -- f
           -- code x65
           "00000000", -- 0
           "00000000", -- 1
           "00000000", -- 2
           "00000000", -- 3
           "00000000", -- 4
           "01111100", -- 5  *****
           "11000110", -- 6 **   **
           "11111110", -- 7 *******
           "11000000", -- 8 **
           "11000000", -- 9 **
           "11000110", -- a **   **
           "01111100", -- b  *****
           "00000000", -- c
           "00000000", -- d
           "00000000", -- e
           "00000000", -- f
           -- code x66
           "00000000", -- 0
           "00000000", -- 1
           "00111000", -- 2   ***
           "01101100", -- 3  ** **
           "01100100", -- 4  **  *
           "01100000", -- 5  **
           "11110000", -- 6 ****
           "01100000", -- 7  **
           "01100000", -- 8  **
           "01100000", -- 9  **
           "01100000", -- a  **
           "11110000", -- b ****
           "00000000", -- c
           "00000000", -- d
           "00000000", -- e
           "00000000", -- f
           -- code x67
           "00000000", -- 0
           "00000000", -- 1
           "00000000", -- 2
           "00000000", -- 3
           "00000000", -- 4
           "01110110", -- 5  *** **
           "11001100", -- 6 **  **
           "11001100", -- 7 **  **
           "11001100", -- 8 **  **
           "11001100", -- 9 **  **
           "11001100", -- a **  **
           "01111100", -- b  *****
           "00001100", -- c     **
           "11001100", -- d **  **
           "01111000", -- e  ****
           "00000000", -- f
           -- code x68
           "00000000", -- 0
           "00000000", -- 1
           "11100000", -- 2 ***
           "01100000", -- 3  **
           "01100000", -- 4  **
           "01101100", -- 5  ** **
           "01110110", -- 6  *** **
           "01100110", -- 7  **  **
           "01100110", -- 8  **  **
           "01100110", -- 9  **  **
           "01100110", -- a  **  **
           "11100110", -- b ***  **
           "00000000", -- c
           "00000000", -- d
           "00000000", -- e
           "00000000", -- f
           -- code x69
           "00000000", -- 0
           "00000000", -- 1
           "00011000", -- 2    **
           "00011000", -- 3    **
           "00000000", -- 4
           "00111000", -- 5   ***
           "00011000", -- 6    **
           "00011000", -- 7    **
           "00011000", -- 8    **
           "00011000", -- 9    **
           "00011000", -- a    **
           "00111100", -- b   ****
           "00000000", -- c
           "00000000", -- d
           "00000000", -- e
           "00000000", -- f
           -- code x6a
           "00000000", -- 0
           "00000000", -- 1
           "00000110", -- 2      **
           "00000110", -- 3      **
           "00000000", -- 4
           "00001110", -- 5     ***
           "00000110", -- 6      **
           "00000110", -- 7      **
           "00000110", -- 8      **
           "00000110", -- 9      **
           "00000110", -- a      **
           "00000110", -- b      **
           "01100110", -- c  **  **
           "01100110", -- d  **  **
           "00111100", -- e   ****
           "00000000", -- f
           -- code x6b
           "00000000", -- 0
           "00000000", -- 1
           "11100000", -- 2 ***
           "01100000", -- 3  **
           "01100000", -- 4  **
           "01100110", -- 5  **  **
           "01101100", -- 6  ** **
           "01111000", -- 7  ****
           "01111000", -- 8  ****
           "01101100", -- 9  ** **
           "01100110", -- a  **  **
           "11100110", -- b ***  **
           "00000000", -- c
           "00000000", -- d
           "00000000", -- e
           "00000000", -- f
           -- code x6c
           "00000000", -- 0
           "00000000", -- 1
           "00111000", -- 2   ***
           "00011000", -- 3    **
           "00011000", -- 4    **
           "00011000", -- 5    **
           "00011000", -- 6    **
           "00011000", -- 7    **
           "00011000", -- 8    **
           "00011000", -- 9    **
           "00011000", -- a    **
           "00111100", -- b   ****
           "00000000", -- c
           "00000000", -- d
           "00000000", -- e
           "00000000", -- f
           -- code x6d
           "00000000", -- 0
           "00000000", -- 1
           "00000000", -- 2
           "00000000", -- 3
           "00000000", -- 4
           "11100110", -- 5 ***  **
           "11111111", -- 6 ********
           "11011011", -- 7 ** ** **
           "11011011", -- 8 ** ** **
           "11011011", -- 9 ** ** **
           "11011011", -- a ** ** **
           "11011011", -- b ** ** **
           "00000000", -- c
           "00000000", -- d
           "00000000", -- e
           "00000000", -- f
           -- code x6e
           "00000000", -- 0
           "00000000", -- 1
           "00000000", -- 2
           "00000000", -- 3
           "00000000", -- 4
           "11011100", -- 5 ** ***
           "01100110", -- 6  **  **
           "01100110", -- 7  **  **
           "01100110", -- 8  **  **
           "01100110", -- 9  **  **
           "01100110", -- a  **  **
           "01100110", -- b  **  **
           "00000000", -- c
           "00000000", -- d
           "00000000", -- e
           "00000000", -- f
           -- code x6f
           "00000000", -- 0
           "00000000", -- 1
           "00000000", -- 2
           "00000000", -- 3
           "00000000", -- 4
           "01111100", -- 5  *****
           "11000110", -- 6 **   **
           "11000110", -- 7 **   **
           "11000110", -- 8 **   **
           "11000110", -- 9 **   **
           "11000110", -- a **   **
           "01111100", -- b  *****
           "00000000", -- c
           "00000000", -- d
           "00000000", -- e
           "00000000", -- f
           -- code x70
           "00000000", -- 0
           "00000000", -- 1
           "00000000", -- 2
           "00000000", -- 3
           "00000000", -- 4
           "11011100", -- 5 ** ***
           "01100110", -- 6  **  **
           "01100110", -- 7  **  **
           "01100110", -- 8  **  **
           "01100110", -- 9  **  **
           "01100110", -- a  **  **
           "01111100", -- b  *****
           "01100000", -- c  **
           "01100000", -- d  **
           "11110000", -- e ****
           "00000000", -- f
           -- code x71
           "00000000", -- 0
           "00000000", -- 1
           "00000000", -- 2
           "00000000", -- 3
           "00000000", -- 4
           "01110110", -- 5  *** **
           "11001100", -- 6 **  **
           "11001100", -- 7 **  **
           "11001100", -- 8 **  **
           "11001100", -- 9 **  **
           "11001100", -- a **  **
           "01111100", -- b  *****
           "00001100", -- c     **
           "00001100", -- d     **
           "00011110", -- e    ****
           "00000000", -- f
           -- code x72
           "00000000", -- 0
           "00000000", -- 1
           "00000000", -- 2
           "00000000", -- 3
           "00000000", -- 4
           "11011100", -- 5 ** ***
           "01110110", -- 6  *** **
           "01100110", -- 7  **  **
           "01100000", -- 8  **
           "01100000", -- 9  **
           "01100000", -- a  **
           "11110000", -- b ****
           "00000000", -- c
           "00000000", -- d
           "00000000", -- e
           "00000000", -- f
           -- code x73
           "00000000", -- 0
           "00000000", -- 1
           "00000000", -- 2
           "00000000", -- 3
           "00000000", -- 4
           "01111100", -- 5  *****
           "11000110", -- 6 **   **
           "01100000", -- 7  **
           "00111000", -- 8   ***
           "00001100", -- 9     **
           "11000110", -- a **   **
           "01111100", -- b  *****
           "00000000", -- c
           "00000000", -- d
           "00000000", -- e
           "00000000", -- f
           -- code x74
           "00000000", -- 0
           "00000000", -- 1
           "00010000", -- 2    *
           "00110000", -- 3   **
           "00110000", -- 4   **
           "11111100", -- 5 ******
           "00110000", -- 6   **
           "00110000", -- 7   **
           "00110000", -- 8   **
           "00110000", -- 9   **
           "00110110", -- a   ** **
           "00011100", -- b    ***
           "00000000", -- c
           "00000000", -- d
           "00000000", -- e
           "00000000", -- f
           -- code x75
           "00000000", -- 0
           "00000000", -- 1
           "00000000", -- 2
           "00000000", -- 3
           "00000000", -- 4
           "11001100", -- 5 **  **
           "11001100", -- 6 **  **
           "11001100", -- 7 **  **
           "11001100", -- 8 **  **
           "11001100", -- 9 **  **
           "11001100", -- a **  **
           "01110110", -- b  *** **
           "00000000", -- c
           "00000000", -- d
           "00000000", -- e
           "00000000", -- f
           -- code x76
           "00000000", -- 0
           "00000000", -- 1
           "00000000", -- 2
           "00000000", -- 3
           "00000000", -- 4
           "11000011", -- 5 **    **
           "11000011", -- 6 **    **
           "11000011", -- 7 **    **
           "11000011", -- 8 **    **
           "01100110", -- 9  **  **
           "00111100", -- a   ****
           "00011000", -- b    **
           "00000000", -- c
           "00000000", -- d
           "00000000", -- e
           "00000000", -- f
           -- code x77
           "00000000", -- 0
           "00000000", -- 1
           "00000000", -- 2
           "00000000", -- 3
           "00000000", -- 4
           "11000011", -- 5 **    **
           "11000011", -- 6 **    **
           "11000011", -- 7 **    **
           "11011011", -- 8 ** ** **
           "11011011", -- 9 ** ** **
           "11111111", -- a ********
           "01100110", -- b  **  **
           "00000000", -- c
           "00000000", -- d
           "00000000", -- e
           "00000000", -- f
           -- code x78
           "00000000", -- 0
           "00000000", -- 1
           "00000000", -- 2
           "00000000", -- 3
           "00000000", -- 4
           "11000011", -- 5 **    **
           "01100110", -- 6  **  **
           "00111100", -- 7   ****
           "00011000", -- 8    **
           "00111100", -- 9   ****
           "01100110", -- a  **  **
           "11000011", -- b **    **
           "00000000", -- c
           "00000000", -- d
           "00000000", -- e
           "00000000", -- f
           -- code x79
           "00000000", -- 0
           "00000000", -- 1
           "00000000", -- 2
           "00000000", -- 3
           "00000000", -- 4
           "11000110", -- 5 **   **
           "11000110", -- 6 **   **
           "11000110", -- 7 **   **
           "11000110", -- 8 **   **
           "11000110", -- 9 **   **
           "11000110", -- a **   **
           "01111110", -- b  ******
           "00000110", -- c      **
           "00001100", -- d     **
           "11111000", -- e *****
           "00000000", -- f
           -- code x7a
           "00000000", -- 0
           "00000000", -- 1
           "00000000", -- 2
           "00000000", -- 3
           "00000000", -- 4
           "11111110", -- 5 *******
           "11001100", -- 6 **  **
           "00011000", -- 7    **
           "00110000", -- 8   **
           "01100000", -- 9  **
           "11000110", -- a **   **
           "11111110", -- b *******
           "00000000", -- c
           "00000000", -- d
           "00000000", -- e
           "00000000", -- f
           -- code x7b {
           "00000000", -- 0
           "00000000", -- 1
           "00001110", -- 2     ***
           "00011000", -- 3    **
           "00011000", -- 4    **
           "00011000", -- 5    **
           "01110000", -- 6  ***
           "00011000", -- 7    **
           "00011000", -- 8    **
           "00011000", -- 9    **
           "00011000", -- a    **
           "00001110", -- b     ***
           "00000000", -- c
           "00000000", -- d
           "00000000", -- e
           "00000000", -- f
           -- code x7c |
           "00000000", -- 0
           "00000000", -- 1
           "00011000", -- 2    **
           "00011000", -- 3    **
           "00011000", -- 4    **
           "00011000", -- 5    **
           "00000000", -- 6
           "00011000", -- 7    **
           "00011000", -- 8    **
           "00011000", -- 9    **
           "00011000", -- a    **
           "00011000", -- b    **
           "00000000", -- c
           "00000000", -- d
           "00000000", -- e
           "00000000", -- f
           -- code x7d }
           "00000000", -- 0
           "00000000", -- 1
           "01110000", -- 2  ***
           "00011000", -- 3    **
           "00011000", -- 4    **
           "00011000", -- 5    **
           "00001110", -- 6     ***
           "00011000", -- 7    **
           "00011000", -- 8    **
           "00011000", -- 9    **
           "00011000", -- a    **
           "01110000", -- b  ***
           "00000000", -- c
           "00000000", -- d
           "00000000", -- e
           "00000000", -- f
           -- code x7e ~
           "00000000", -- 0
           "00000000", -- 1
           "01110110", -- 2  *** **
           "11011100", -- 3 ** ***
           "00000000", -- 4
           "00000000", -- 5
           "00000000", -- 6
           "00000000", -- 7
           "00000000", -- 8
           "00000000", -- 9
           "00000000", -- a
           "00000000", -- b
           "00000000", -- c
           "00000000", -- d
           "00000000", -- e
           "00000000", -- f
           -- code x7f
           "00000000", -- 0
           "00000000", -- 1
           "00000000", -- 2
           "00000000", -- 3
           "00010000", -- 4    *
           "00111000", -- 5   ***
           "01101100", -- 6  ** **
           "11000110", -- 7 **   **
           "11000110", -- 8 **   **
           "11000110", -- 9 **   **
           "11111110", -- a *******
           "00000000", -- b
           "00000000", -- c
           "00000000", -- d
           "00000000", -- e
           "00000000"  -- f
           );
        begin
            --return X <= 8 and Y <= 16 and ROM((char * 16) + Y)(9 - X) = '1';
            return ROM((CHARACTER'POS(char) * 16) + Y)(9 - X) = '1';
        end draw_char;
        

--        The MIT License (MIT)
        
--        Copyright (c) 2016 Dries007
        
--        Permission is hereby granted, free of charge, to any person obtaining a copy
--        of this software and associated documentation files (the "Software"), to deal
--        in the Software without restriction, including without limitation the rights
--        to use, copy, modify, merge, publish, distribute, sublicense, and/or sell
--        copies of the Software, and to permit persons to whom the Software is
--        furnished to do so, subject to the following conditions:
        
--        The above copyright notice and this permission notice shall be included in all
--        copies or substantial portions of the Software.
        
--        THE SOFTWARE IS PROVIDED "AS IS", WITHOUT WARRANTY OF ANY KIND, EXPRESS OR
--        IMPLIED, INCLUDING BUT NOT LIMITED TO THE WARRANTIES OF MERCHANTABILITY,
--        FITNESS FOR A PARTICULAR PURPOSE AND NONINFRINGEMENT. IN NO EVENT SHALL THE
--        AUTHORS OR COPYRIGHT HOLDERS BE LIABLE FOR ANY CLAIM, DAMAGES OR OTHER
--        LIABILITY, WHETHER IN AN ACTION OF CONTRACT, TORT OR OTHERWISE, ARISING FROM,
--        OUT OF OR IN CONNECTION WITH THE SOFTWARE OR THE USE OR OTHER DEALINGS IN THE
--        SOFTWARE.
 
        function draw_string(scanX : natural; scanY : natural; posX : natural; posY : natural; s : string; center : boolean; size : natural) return boolean is
            constant charW : natural := 8 * size;
            constant charWsp : natural := charW + 2;
            constant charH : natural := 16 * size;
            constant width : natural := charWsp * s'LENGTH;
            constant height : natural := charH;
            variable x : natural := posX;
            variable y : natural := posY;
            variable char : natural;
            variable subX : natural;
            begin
                if (center) then
                    x := x - (width / 2);
                    y := y - (height / 2);
                end if;
            
                if (scanX < x or scanY < y) then
                    return false;
                end if;
                
                if (scanX - x > width or scanY - y > height) then
                    return false;
                end if;
                
                x := scanX - x;
                y := scanY - y;
                
                subX := x mod charWsp;
                char := (x / charWsp) + 1;
                
                return draw_char(subX / size, y / size, s(char));
        end draw_string;
begin
	VGA: entity work.vga
        port map (
            CLK_I => clk,
            VGA_RED_O => vgaRed,
            VGA_BLUE_O => vgaBlue,
            VGA_GREEN_O => vgaGreen,
            VGA_HS_O => Hsync,
            VGA_VS_O => Vsync,
            X => X,
            Y => Y,
            R => Red,
            G => Green,
            B => Blue
        );
    
--	DB_U: entity work.debounce
--			port map (
--				clk => clk,
--				button => btnU,
--				result => btnU_DB
--			);

--	DB_D: entity work.debounce
--			port map (
--				clk => clk,
--				button => btnD,
--				result => btnD_DB
--			);
    	
	sevenSegDisplay : Sequential_7Segments_Decoder
	       port map (
	            clk => clk,
	            value(3 downto 0) => in0,
	            value(7 downto 4) => in1,
	            value(11 downto 8)=> in2,
	            value(15 downto 12)=> in3,
	            segs => seg,
	            dp => dp,
	            channels => an,
	            RESET => '0'   
	       );
	       
	 PS2Key : ps2keyboard
	       port map(
	                  resetn => '1', 
	                  clock => clk,
                      ps2c => ps2c_in, 
                      ps2d => ps2d_in,
                      DOUT => Dout,
                      code => code_out
                              );
                              
	--Setting the motion up or down
        process(reset, Dout)
        begin
        
                        if( reset = '1' ) then --Resetting the game
                            moveUp <= '0';
                            moveDown <= '0';              
                        else
                            --Direction
                            if( Dout(7 downto 0) = "01110101") then
                                moveUp <= '1';
                                moveDown <= '0';
                            elsif( Dout(7 downto 0) = "01110010") then
                                moveUp <= '0';
                                moveDown <= '1';
                            end if;
                        end if;
                    
                end process;
    
    --Motion
    process( clk, reset, moveUp, moveDown)
    begin
         if( rising_edge(clk) ) then
            clk_cnt <= clk_cnt + 1;
            if( reset = '1' ) then
                posX <= centerX;
                posY <= centerY;
                gameOver <= '0';
            elsif( clk_cnt >= 500000) then
                clk_cnt <= 0;
                
                if( gameOver = '0' ) then --For less energy use
                    --Motion
                    if( moveUp = '1' and posY >= speedOfGuy) then
                         posY <= posY - speedOfGuy;
                    elsif( moveDown = '1' and posY <= 1024 - sizeOfGuy + speedOfGuy) then
                        posY <= posY + speedOfGuy;
                    end if; 
                    
                    --Collision
                    if( ( posY + sizeOfGuy >= currentUpEdge and posY <= currentUpEdge + heightOfBar)
                          or ( posY + sizeOfGuy >= currentDownEdge and posY <= currentDownEdge + heightOfBar)
                          or posY <= speedOfGuy or posY >= 1024 - sizeOfGuy ) then
                        gameOver <= '1';
                    end if; 
                end if;
                     
            end if;
         end if;
    end process;
    
	--Mechanics for the motion of bars
	process( clk )    
	begin
	   if (rising_edge(clk)) then
           frame_count <= frame_count + 1;
           if( reset = '1') then --Resetting the game
               indexUpBarNext <= 0;
               upBarXPositions <= (1280, 1280 + upBarLengths(0), 1280 + upBarLengths(0) + upBarLengths(1),
                                   1280 + upBarLengths(0) + upBarLengths(1) + upBarLengths(2),
                                   1280 + upBarLengths(0) + upBarLengths(1) + upBarLengths(2) + upBarLengths(3) );
               upBarYPositions <= (350,300,250,200,250);
               upBarLengths <= ( 256,256, 256, 256,256);
               
               indexDownBarNext <= 0;
               downBarXPositions <= (centerX, centerX + downBarLengths(0), centerX + downBarLengths(0) + downBarLengths(1),
                                     centerX + downBarLengths(0) + downBarLengths(1) + downBarLengths(2),
                                     centerX + downBarLengths(0) + downBarLengths(1) + downBarLengths(2) + downBarLengths(3) );
               downBarYPositions <= (700, 580, 610, 640,640);
               downBarLengths <= ( 256,256,256,256,256);
           elsif (frame_count >= 500000) then
               frame_count <= 0;
               if( gameOver = '0' ) then
                   for i in 0 to 4 loop
                      upBarXPositions(i) <= upBarXPositions(i) - speedOfBars;
                      downBarXPositions(i) <= downBarXPositions(i) - speedOfBars;
                      if( upBarXPositions(i) + upBarLengths(i) <= 0) then
                          --Up Bars
                          upBarXPositions(i) <= 1280;
                          upBarLengths(i) <= upBarLengthsNext( indexUpBarNext);
                          upBarYPositions(i) <= upBarYPositionsNext( indexUpBarNext);
                          if( indexUpBarNext >= 99) then
                               indexUpBarNext <= 0;
                          else
                               indexUpBarNext <= indexUpBarNext + 1;
                          end if;
                       end if;
                           
                       if ( downBarXPositions(i) + downBarLengths(i) <= 0) then
                         --Down Bars
                         downBarXPositions(i) <= 1280;
                         downBarLengths(i) <= downBarLengthsNext( indexDownBarNext);
                         downBarYPositions(i) <= downBarYPositionsNext( indexDownBarNext);
                         if( indexDownBarNext >= 99) then
                             indexDownBarNext <= 0;
                         else
                             indexDownBarNext <= indexDownBarNext + 1;
                         end if;
                         
                      end if;
                    end loop;
               end if;
               
           end if;
       end if;
	end process;
	
	--Mechanis for current edge of up bar, no need to divide clk or clk in sensivity list since upBarXPositions change
	-- with the rate of the frame
	process( clk, upBarXPositions, posX, gameOver, upBarLengths, upBarYPositions)
	begin
	   if (rising_edge(clk)) then
	       curUp_cnt <= curUp_cnt + 1;
	       if( reset = '1') then
	           curUp_cnt <= 0;
	       elsif( curUp_cnt >= 900) then
	           curUp_cnt <= 0;
	           if( gameOver = '0' ) then
                  for i in 0 to 4 loop
                     if( posX + sizeOfGuy >= upBarXPositions(i)  and posX <= upBarXPositions(i) + upBarLengths(i) - sizeOfGuy ) then
                         currentUpEdge <= upBarYPositions(i);
                         exit;
                     else
                         currentUpEdge <= 0;    
                     end if;
                  end loop;
              end if; 
	       end if;
	   end if; 
	end process;
	
	--Mechanis for current edge of down bar, no need to divide clk or clk in sensivity list since upBarXPositions change
    -- with the rate of the frame
	process( clk, downBarXPositions, posX, gameOVer, downBarLengths, downBarYPositions)
    begin
        if( rising_edge(clk) ) then
            curDown_cnt <= curDown_cnt + 1;
            if( reset = '1') then
                curDown_cnt <= 0;
            elsif( curDown_cnt >= 900) then
                curDown_cnt <= 0;
                if( gameOver = '0' ) then
                    for i in 0 to 4 loop
                       if( posX + sizeOfGuy >= downBarXPositions(i)  and posX <= downBarXPositions(i) + downBarLengths(i) - sizeOfGuy ) then
                           currentDownEdge <= downBarYPositions(i);
                           exit;
                       else
                           currentDownEdge <= 1024;    
                       end if;
                   end loop;
                end if; 
            end if;
        end if;
    end process;
	
	--Timer for score
	process( clk)
	begin
        if( rising_edge(clk)) then
            score_cnt <= score_cnt + 1;
            if( reset = '1') then
                score_cnt <= 0;
                score <= 0;
            elsif( score_cnt >= 10000000) then
                score_cnt <= 0;
                if( gameOver = '0' ) then
                    score <= score + 1;
                end if;
            end if;
        end if;
	end process;
	
	--Showing the socre on 7 segment display
	process( score)
	variable integer0: natural range 0 to 9;
	variable integer1: natural range 0 to 9;
	variable integer1mod: natural range 0 to 99;
	variable integer2: natural range 0 to 9;
	variable integer2mod: natural range 0 to 999;
	variable integer3: natural range 0 to 9;
	begin
	   integer0 := score mod 10;
	   in0 <=  conv_std_logic_vector(integer0,4);
	   
	   integer1mod := score mod 100;
	   integer1 := integer1Mod / 10;
	   in1 <= conv_std_logic_vector(integer1,4);
	   
	   integer2mod := score mod 1000;
	   integer2 := integer2mod / 100;
	   in2 <= conv_std_logic_vector(integer2,4);
	   
	   integer3 := score / 1000;
	   in3 <= conv_std_logic_vector(integer3,4);
	end process;
	
	--Adjusting the speed according to score
	process( clk, speed_sw)
	begin
	   if( rising_edge(clk) ) then
	      if( reset = '1' ) then
              speedOfGuy <= 1;
              speedOfBars <= 1;
          elsif ( speed_sw = "000") then --000
              speedOfGuy <= 1;
              speedOfBars <= 1;
          elsif( speed_sw  = "001") then --001
              speedOfGuy <= 2;
              speedOfBars <= 2;
          elsif( speed_sw  = "010") then --010
              speedOfGuy <= 3;
              speedOfBars <= 3;
          elsif( speed_sw  = "011") then --011
              speedOfGuy <= 4;
              speedOfBars <= 4;
          else
            speedOfBars <=5;
          
          end if;
	   end if;
	end process;
	
	--Drawing the video
	process( X, Y, gameOver, posX, posY, upBarXPositions, upBarYPositions, upBarLengths, downBarYPositions, downBarXPositions, downBarLengths)
	begin
	    if( gameOver = '1' ) then
	       if (draw_string(X, Y, centerX, centerY, "GAME OVER!", true, 5)) then
	           Red <= 15;
               Green <= 15;
               Blue <= 0;
	       else
	           Red <= 0;
	           Green <= 0;
	           Blue <= 0;
	       end if;
	    else
	       --Guy
            if( Y > posY and Y < posY + sizeOfGuy and X > posX and X < posX + sizeOfGuy ) then
                    if( gameOver = '1') then
                    Red <= 15;
                    Green <= 15;
                    Blue <= 0;
                    else
                    Red <= 15;
                    Green <= 0;
                    Blue <= 0;
                    end if;

--            else        
--            --Bars
--            for I in 0 to 3 loop -- Not working for some reasons which might be timing issues or if/else structure
--                  if( Y > upBarYPositions(i) - heightOfBar/2 and Y < upBarYPositions(i) + heightOfBar/2
--                           --and  X > barPosX - lengthOfBar/2 + I*lengthOfBar
--                           --and X < barPosX + lengthOfBar/2 + I*lengthOfBar ) then
--                           ) then 
--                    Red <= 0;
--                    Green <= 15;
--                    Blue <= 0;
                    
--                    else
--                    Red <= 0;
--                    Green <= 0;
--                    Blue <= 0;
--                  end if;
--            end loop;

            --Bars
            --Up Bars
            elsif( Y > upBarYPositions(0) and Y < upBarYPositions(0) + heightOfBar
                                   and  X > upBarXPositions(0)
                                   and X < upBarXPositions(0) + upBarLengths(0)) then
                Red <= 0;
                Green <= 15;
                Blue <= 0;
            elsif( Y > upBarYPositions(1) and Y < upBarYPositions(1) + heightOfBar
                                   and  X > upBarXPositions(1)
                                   and X < upBarXPositions(1) + upBarLengths(1) ) then
                Red <= 0;
                Green <= 15;
                Blue <= 0;
                            
            elsif( Y > upBarYPositions(2) and Y < upBarYPositions(2) + heightOfBar
                                   and  X > upBarXPositions(2) 
                                   and X < upBarXPositions(2) + upBarLengths(2) ) then
                Red <= 0;
                Green <= 15;
                Blue <= 0;
                                        
            elsif( Y > upBarYPositions(3) and Y < upBarYPositions(3) + heightOfBar
                                   and  X > upBarXPositions(3)
                                   and X < upBarXPositions(3) + upBarLengths(3) ) then
                Red <= 0;
                Green <= 15;
                Blue <= 0;
            elsif( Y > upBarYPositions(4) and Y < upBarYPositions(4) + heightOfBar
                                   and  X > upBarXPositions(4)
                                   and X < upBarXPositions(4) + upBarLengths(4) ) then
                Red <= 0;
                Green <= 15;
                Blue <= 0;
            
            elsif( Y > downBarYPositions(0) and Y < downBarYPositions(0) + heightOfBar
                                   and  X > downBarXPositions(0)
                                   and X < downBarXPositions(0) + downBarLengths(0)) then
                Red <= 0;
                Green <= 0;
                Blue <= 15;
            elsif( Y > downBarYPositions(1) and Y < downBarYPositions(1) + heightOfBar
                                   and  X > downBarXPositions(1)
                                   and X < downBarXPositions(1) + downBarLengths(1) ) then
                Red <= 0;
                Green <= 0;
                Blue <= 15;
                            
            elsif( Y > downBarYPositions(2) and Y < downBarYPositions(2) + heightOfBar
                                   and  X > downBarXPositions(2) 
                                   and X < downBarXPositions(2) + downBarLengths(2) ) then
                Red <= 0;
                Green <= 0;
                Blue <= 15;
                                        
            elsif( Y > downBarYPositions(3) and Y < downBarYPositions(3) + heightOfBar
                                   and  X > downBarXPositions(3)
                                   and X < downBarXPositions(3) + downBarLengths(3) ) then
                Red <= 0;
                Green <= 0;
                Blue <= 15;
            elsif( Y > downBarYPositions(4) and Y < downBarYPositions(4) + heightOfBar
                                   and  X > downBarXPositions(4)
                                   and X < downBarXPositions(4) + downBarLengths(4) ) then
                Red <= 0;
                Green <= 0;
                Blue <= 15;
                
            --Background
            else
               Red <= 0;
               Green <= 0;
               Blue <= 0;         
            end if;
	    end if;

	end process;
end Behavioral;